module Firmware (
	input clk

 
);

endmodule